version https://git-lfs.github.com/spec/v1
oid sha256:53ed3ef12f0cb34aa427a91a0b5e885b3aa4d9d800738e1111b2b2ed188ed140
size 2411
