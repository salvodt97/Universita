version https://git-lfs.github.com/spec/v1
oid sha256:7cf529f74e029741213b1e69d8dc6e7fad3c3baa89e37977ed39cfd204144dab
size 326
