version https://git-lfs.github.com/spec/v1
oid sha256:5597dc377f906bff34951756cc64c0570adfed31a19fb3eb0b6d649a4599952d
size 3273
