version https://git-lfs.github.com/spec/v1
oid sha256:f9cdc0332020b29278bb8666bb844070e17e6721137a2ade0debe5381d338378
size 277
