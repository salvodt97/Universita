version https://git-lfs.github.com/spec/v1
oid sha256:ec5575833e68e01a2101d6ea0a153afa83d48904df04c85c3de6cb01744a3800
size 1997
