version https://git-lfs.github.com/spec/v1
oid sha256:0a3adb154ee130e77b6d6589a629b23ae161eb650d0aa5532ce322a7f0330aaa
size 2021
