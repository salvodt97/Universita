version https://git-lfs.github.com/spec/v1
oid sha256:a8a26b907915eef4f7385f874c89b0c6daca1adef8f9aba3c524d84c2878abbe
size 2677
