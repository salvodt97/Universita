version https://git-lfs.github.com/spec/v1
oid sha256:3c1aba8946c38ba2b7499e8359eb4f6f188527190337a332b9a90ad4ede4e41b
size 709
