version https://git-lfs.github.com/spec/v1
oid sha256:0af10567998195852c22a8c220abb3b7fb58ce90231b722553939556417b53a3
size 636
