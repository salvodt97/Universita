version https://git-lfs.github.com/spec/v1
oid sha256:299060a15620d43be3c49d19689a7cb4fc1a2b84ad027bb68b04c56520fb078a
size 1172
