version https://git-lfs.github.com/spec/v1
oid sha256:0533646f45cccf926cb46a5496953525cc6c75f50eaa4402f4f1447a88c46083
size 983
