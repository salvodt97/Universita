version https://git-lfs.github.com/spec/v1
oid sha256:90d2a14d5b13f1207dcafc1f95e08181a130e1780a29d5f61de5e771d959fcf2
size 1120
