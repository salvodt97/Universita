version https://git-lfs.github.com/spec/v1
oid sha256:236c97a3d223c186015b0d383447dedfb177e9c697bf585e5d61709ccdd5872f
size 773
