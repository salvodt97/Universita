version https://git-lfs.github.com/spec/v1
oid sha256:acfee049f3014e60ca56044a4d3cc4a694c6d53120c1a660064a893806651e47
size 1218
