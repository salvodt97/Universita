version https://git-lfs.github.com/spec/v1
oid sha256:b5657b10819ecc86c4c3e06a540d194598a00bc4063f6a584a98f0bae646890d
size 668
