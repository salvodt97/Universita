version https://git-lfs.github.com/spec/v1
oid sha256:972b99de65b7c07304df06294f6d2bcaa1b422f0e35e41cb917ef53e395579ee
size 5954
