version https://git-lfs.github.com/spec/v1
oid sha256:eccde8f2ace052f92d65244283e7bf389b9a728bccb2a82332b299d39fe5fea6
size 999
