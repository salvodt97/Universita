version https://git-lfs.github.com/spec/v1
oid sha256:11d4fd571ea97c1ba10d595bed4136a2cd5733bd69e58849400b99d982e2214a
size 845
