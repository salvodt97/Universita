version https://git-lfs.github.com/spec/v1
oid sha256:a0c20970d3a403e54ef9b90a31037a6dc487c0abaf40aefc34dc69ad05d6dad6
size 2547
