version https://git-lfs.github.com/spec/v1
oid sha256:aa95d702cfd8f72dbe42918e6577430d33b6bc4fe9c4f0d9659639cf8941cfe6
size 1191
