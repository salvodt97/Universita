version https://git-lfs.github.com/spec/v1
oid sha256:a6d16ba7de936109088c881eedcf3031c26c006ac596fe75b1babda39fcbe0a0
size 774
