version https://git-lfs.github.com/spec/v1
oid sha256:6ce19d200730d235e5cd561c75d525c5666415c348f3da3fb848fafdcd4b3a3d
size 1570
