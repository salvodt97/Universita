version https://git-lfs.github.com/spec/v1
oid sha256:2b074f8e802a176c20a3a9e51d8c82ee14cec336a02667288f991f318b351565
size 3068
