version https://git-lfs.github.com/spec/v1
oid sha256:077ce82c15514e7c78e067338bf2beeb5b0d68db4f66e41d098301224e048a33
size 879
