version https://git-lfs.github.com/spec/v1
oid sha256:e5de74faa0c5b22b2521221e4e233d3f0dace8693100072474e1dac0145f0518
size 1987
