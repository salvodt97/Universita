version https://git-lfs.github.com/spec/v1
oid sha256:ad3b8b91ece2e6d44dd70633b9c53585bca50f10255ddeb1bf26364ff29ede07
size 432
