version https://git-lfs.github.com/spec/v1
oid sha256:238a3487e43bd60eb63f3d1f12cec65f40fe418a362ced55e0537d43c17af480
size 3016
