version https://git-lfs.github.com/spec/v1
oid sha256:390985bcc39faea767ebc0455aef0ed192911752d826f682976a793d485f807f
size 1010
