version https://git-lfs.github.com/spec/v1
oid sha256:f5cf3d13f00596deed42b8077a55fa614425a426e5cc7e60fc490288c84f61d8
size 275
