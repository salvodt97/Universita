version https://git-lfs.github.com/spec/v1
oid sha256:88d523835d97a166d375ae15b7f9dd5e475af6f3579bb505fdb56d611b892c1f
size 2068
