version https://git-lfs.github.com/spec/v1
oid sha256:b29465f5fef08f2f38dde15fb1ce296dca56a7c59ff6401e7eaeb13eef780356
size 1569
