version https://git-lfs.github.com/spec/v1
oid sha256:a95f7d4a63f219cbb643c8a8b2f305a1f9ba038a6b88022db3f241712ad2426f
size 2375
