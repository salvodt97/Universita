version https://git-lfs.github.com/spec/v1
oid sha256:46b2adb5fcceaef49ec2cef86e26b48a95478039aeb55d955f49cf189a602878
size 8836
