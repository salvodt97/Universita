version https://git-lfs.github.com/spec/v1
oid sha256:18e27c0e49fc71c585def2a4c90dc8a8db220fbb30c6a350d1f033cc406f78e6
size 600
