version https://git-lfs.github.com/spec/v1
oid sha256:aefa526fc2fe2a66bfdbce23442358df916d4775192f4c5049bc2964e1338b54
size 1837
