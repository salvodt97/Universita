version https://git-lfs.github.com/spec/v1
oid sha256:ad3d5e7a2c1881c885fb87182c2a49d639c4f149210533bad99d60d89ca2a339
size 972
