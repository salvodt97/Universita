version https://git-lfs.github.com/spec/v1
oid sha256:706453fa69b48a0606e6f840e33ca290bbdfd47abcb36be371303edeb82391ab
size 1279
