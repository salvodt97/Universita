version https://git-lfs.github.com/spec/v1
oid sha256:46fbab8df2b3208473ff3ecf69ab328df59550dc4eec59f52299fea31ece54aa
size 673
