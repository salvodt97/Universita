version https://git-lfs.github.com/spec/v1
oid sha256:8db01ebaeffc0e3aeef507a328d4d60cac06d3eacd59fa0c701eb46d18c61c4b
size 1183
