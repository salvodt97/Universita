version https://git-lfs.github.com/spec/v1
oid sha256:58f7ff99803cee0e541d3dc16687d2a2fe05034c4c8b19f8ba8058ff28296d45
size 563
