version https://git-lfs.github.com/spec/v1
oid sha256:13eaaacfbab13bbfc1a63bbb414ab75813da52008b5aa40c5bb2cc92f0637800
size 961
