version https://git-lfs.github.com/spec/v1
oid sha256:3f2b3c5bfb901d2f5f242358613bf069ed0ecb771f821902d38fd29797e6a982
size 1591
