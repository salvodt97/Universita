version https://git-lfs.github.com/spec/v1
oid sha256:cc63d5a71f6c6a04169f186a0520ecb4b0962d774186baabadb0dd68536a50c4
size 28967
