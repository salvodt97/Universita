version https://git-lfs.github.com/spec/v1
oid sha256:2c87f2ece2eb0ad2dcb5b13687a16145304dd7773f5b7d4c12fe3f89887911fb
size 2824
