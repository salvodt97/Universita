version https://git-lfs.github.com/spec/v1
oid sha256:b6e1c1ea95e13d67a011d9e5bc5e17e6dd9b199955c7c130ea38df93d4ba0e60
size 984
