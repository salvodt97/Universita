version https://git-lfs.github.com/spec/v1
oid sha256:aca487359220445cec3cafe1bb20dda265d6c229596e14d50ae7424b0bcb4eef
size 1030
