version https://git-lfs.github.com/spec/v1
oid sha256:1b26c7a39a746145841c0f00d447797fd8882cffc775a1fc4cb58422dfa04de4
size 2136
