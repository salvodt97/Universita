version https://git-lfs.github.com/spec/v1
oid sha256:f742afb44ed19c73ff3688a0c159c2c7585fef3288b0a051778c2cacae68f8db
size 28969
