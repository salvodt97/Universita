version https://git-lfs.github.com/spec/v1
oid sha256:6b992b266e85a86c44350b12791f55b057a5e61a6b4278e00315813c24b420ad
size 796
