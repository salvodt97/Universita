version https://git-lfs.github.com/spec/v1
oid sha256:2bec22d6b49195ebdd3f3e2ece4afd803e205bb4e72973c372c9fa9fa9e11541
size 3232
