version https://git-lfs.github.com/spec/v1
oid sha256:58a24489b7c05bb744d6bc22e717d87baef4086eed6ac4ff368f7334a96033d6
size 591
