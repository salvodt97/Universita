version https://git-lfs.github.com/spec/v1
oid sha256:0e403ed6a83548b6c0b47720f086f58c1ab57c6c9b04adb839bfa8d26508a715
size 671
