version https://git-lfs.github.com/spec/v1
oid sha256:581f6329195fba3f803691c09dceae27804d1582dd31c33b9a5554aa79b1de8b
size 1933
