version https://git-lfs.github.com/spec/v1
oid sha256:290ccaebeba031bfb12582ffe9abc9de0facd86102bb9f701f3818789d9640d4
size 1118
