version https://git-lfs.github.com/spec/v1
oid sha256:2715c88467dacc2e700efb81ab22d153ad8f71692936ee79c96648185bfe34ce
size 1090
