version https://git-lfs.github.com/spec/v1
oid sha256:3ba61ec8bfc36f40fd87b84da9b4939215891462eecc5bf5defd488260f4a0ec
size 825
