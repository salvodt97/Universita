version https://git-lfs.github.com/spec/v1
oid sha256:d9fed7fdf38b728410bc0cf16967999990cc7a098a5d473312de350e6d4a2856
size 1067
