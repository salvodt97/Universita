version https://git-lfs.github.com/spec/v1
oid sha256:f34070a151d39622ceb275bfca65b5bd7e5711e875cb548700a3a509d307019d
size 4097
