version https://git-lfs.github.com/spec/v1
oid sha256:85077510859c45eec8da29d1b873e3f3446ab182065c4b4e4cef15966a8a5dfc
size 548
