version https://git-lfs.github.com/spec/v1
oid sha256:167d35e643c02fa8d0b19355bc7b7a222040c0717aab8a703fe335304e27727c
size 1194
