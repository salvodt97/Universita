version https://git-lfs.github.com/spec/v1
oid sha256:ccd5156d09f91a6de42896300f5523cb692403f6630a0935b3afa9e207d90055
size 700
