version https://git-lfs.github.com/spec/v1
oid sha256:503e7e3a01d3b1654abf7495bea0f5d23f3f9e757a5a101f427ca292351dacdc
size 1189
