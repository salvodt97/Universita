version https://git-lfs.github.com/spec/v1
oid sha256:a7a78305630f93765f987c2bfec0dfca7e48545f314a431064b534dac9b16cd1
size 1917
