version https://git-lfs.github.com/spec/v1
oid sha256:2f7f38913e92883318e8b5159c9d8a2682a92611586e468ae85437b51fdbc9d7
size 541
