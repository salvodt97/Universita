version https://git-lfs.github.com/spec/v1
oid sha256:0ad90e74134b629dec5bff06f25aa357e240641d33a307f8a789992b0d38eb65
size 2056
