version https://git-lfs.github.com/spec/v1
oid sha256:485918788aaefc6b63ad158ee233bf9b22ded9fcce7fc8aa1f2a23fecb44b620
size 1067
