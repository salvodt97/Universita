version https://git-lfs.github.com/spec/v1
oid sha256:896aae18e40f394a3dc5c638f2f958b7aa7475067b15366871e2cac8227d4fb4
size 692
