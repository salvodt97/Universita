version https://git-lfs.github.com/spec/v1
oid sha256:00e5f3e76afd9f13e88a948b5a29624aacfef66f8cf9040398f22a5cce24b13e
size 861
