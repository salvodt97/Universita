version https://git-lfs.github.com/spec/v1
oid sha256:a92130d2c4708b39f6cf4950c34ec139e37ad03e414c5d6e3fb8cbb3a2c6a757
size 2655
