version https://git-lfs.github.com/spec/v1
oid sha256:c7112519aee824fbc64c905300b132529ef0fe4b0f7c96244391aae0c9fa3749
size 1184
