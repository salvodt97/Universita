version https://git-lfs.github.com/spec/v1
oid sha256:ff859c5e6464423d466e47752f933531c46931d1f864b5294424bd8b15b0e04b
size 25737
