version https://git-lfs.github.com/spec/v1
oid sha256:07f3d74235b0a26f70be44298fa9bf4cb8f3a3446d3c67c5dc044ce9e7093157
size 5953
