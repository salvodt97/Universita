version https://git-lfs.github.com/spec/v1
oid sha256:91f80c6ce375af92b132b5468b92504f41324af2d1cbdc0ca827dd1f98ffa3f3
size 2052
