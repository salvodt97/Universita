version https://git-lfs.github.com/spec/v1
oid sha256:449d8d39680a1d5019efb9552e1edc7961d06aff1337c2482ad6f6e2f98c9be0
size 841
