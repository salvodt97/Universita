version https://git-lfs.github.com/spec/v1
oid sha256:487dbf40280770b0116c025f0beb0d83d27d116c8d2ebdd4286b25685824f359
size 861
