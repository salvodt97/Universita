version https://git-lfs.github.com/spec/v1
oid sha256:2cf68411bf3b16c2f94a397ed56f5b15b80349efa7a009c1dbc06af3a3a2025a
size 498
