version https://git-lfs.github.com/spec/v1
oid sha256:c25173ba6c1864e7d39c6a19aafa4fdd841b2d7926db174d08c3629fea3859d8
size 2159
