version https://git-lfs.github.com/spec/v1
oid sha256:d24056a0aa2ec899939634917d9ca78d40b3df0cab2aa8ce841d1a9c41a135f1
size 714
