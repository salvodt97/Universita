version https://git-lfs.github.com/spec/v1
oid sha256:ee8e0032dca58b0c345d683e065e87390c85a28efdaaf19d073071bdbaf141a6
size 1162
