version https://git-lfs.github.com/spec/v1
oid sha256:d1dc318b27caea1a5c0ec70d69c2142dba8bf3601b750390960d20cfdffef2df
size 845
