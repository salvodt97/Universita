version https://git-lfs.github.com/spec/v1
oid sha256:2537d6519d98a22679abe475c8fb73608a0d7f6287b62f01e97966a27fd6d589
size 1916
