version https://git-lfs.github.com/spec/v1
oid sha256:51f50ab6ab5e24b27db538ec44892d7d90ee931295481d7133838b2585e19861
size 1164
