version https://git-lfs.github.com/spec/v1
oid sha256:463b3ecf61646956a985d50bfbd60933147e1f3236c96608387ba168d8107b03
size 472
