version https://git-lfs.github.com/spec/v1
oid sha256:d58a4096497d1ea142c06ba4b80570b3d59730d48d9185c7d8faffb5ff63d854
size 759
