version https://git-lfs.github.com/spec/v1
oid sha256:d8348cecc344980d789fef1c54e1222b90da3af14ae869375c5b72c5408dbca5
size 3456
