version https://git-lfs.github.com/spec/v1
oid sha256:45c603facc71d322ff2d1316ceb67392d0a734188d109f9bd5a4916986e6ea0e
size 964
