version https://git-lfs.github.com/spec/v1
oid sha256:9370669878c012ef97c0bcb121839aff3af5e2fbcc1f29f61566f666115b9a27
size 1406
