version https://git-lfs.github.com/spec/v1
oid sha256:ad4fc5cf64539aabfa3a2bf06afa543818e4c685537ed0a885ff57717eb43ea0
size 719
