version https://git-lfs.github.com/spec/v1
oid sha256:ce4fe7dd524b1dfd8cc5db72dc34a637dfd3b4b35f405a3e8179aa974c27f9a2
size 674
