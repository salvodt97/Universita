version https://git-lfs.github.com/spec/v1
oid sha256:7b2499dcaf3c1e8811d2d70074350b408232d59eee46db1ac35c3e0e9f337f58
size 3041
