version https://git-lfs.github.com/spec/v1
oid sha256:10210d475424c45e6ce98ba919c2b5de77d753cac59e4fc098821609f11506fa
size 869
