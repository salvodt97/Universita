version https://git-lfs.github.com/spec/v1
oid sha256:f4e8ad4e2434cef2da224449da0ae59afe48f16dbf00bf82a8ba196683123bf4
size 799
