version https://git-lfs.github.com/spec/v1
oid sha256:cfb961cd0cd3d13c51719ab027ab094ee4be34464485d1985ef8261efcdc2b2c
size 794
