version https://git-lfs.github.com/spec/v1
oid sha256:82b698e2f4b0ca49da61b00d9ddba9408757ad3db3c611b4a40a51dcdd72ddac
size 272
