version https://git-lfs.github.com/spec/v1
oid sha256:8248238c2dbeea69f0ae3cdef0c915207f5bd263b2430ef315a9fce095c06ceb
size 1809
