version https://git-lfs.github.com/spec/v1
oid sha256:f4b20087a08cc78059142ef5cf04470c8c09984f19b849732594ceabfb9fb64c
size 1017
