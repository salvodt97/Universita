version https://git-lfs.github.com/spec/v1
oid sha256:9a401d41339ea9016324afce0c06a67f246ee33a0c28b7811eaa175ba7ba828e
size 835
