version https://git-lfs.github.com/spec/v1
oid sha256:b64796204ba170abe5754723a87fedce56756db96cdd44f44b63dcb81ce4cbdd
size 1129
