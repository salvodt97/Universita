version https://git-lfs.github.com/spec/v1
oid sha256:d5eed4bb58a4404016cd51ddcc3207a80142c8c7d0c5d33d66e778a194ca0ce1
size 1805
