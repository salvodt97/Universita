version https://git-lfs.github.com/spec/v1
oid sha256:32f392277c6c0fc4479754146a9cd7f2a944afc112b5e7753fe1684a5b527d46
size 3109
