version https://git-lfs.github.com/spec/v1
oid sha256:5e1f9613c5186efb5423f87573ab516f8e2c9e7ff8c62b4cca85b5cecf3dce6c
size 506
