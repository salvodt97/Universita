version https://git-lfs.github.com/spec/v1
oid sha256:e122958a5115166d08bf99c2a66bf37f0d8f384f32b2d55ccbdc6d2ea8be7e8b
size 949
