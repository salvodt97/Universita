version https://git-lfs.github.com/spec/v1
oid sha256:90851fdcdf9048d74ebf1f7f9ea5b893ef277a2944108842a0241ee93b10fe8c
size 4308
