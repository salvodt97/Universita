version https://git-lfs.github.com/spec/v1
oid sha256:9c0af472cfe3221590aeac749341b4e14887490c9bbdda1c6a5c56a8095dbbaf
size 4116
