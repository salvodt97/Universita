version https://git-lfs.github.com/spec/v1
oid sha256:190370ad4ffff10ff766fd1a3786ed50236aec52a7bc5766851feb23b6987ec5
size 867
