version https://git-lfs.github.com/spec/v1
oid sha256:ab38fe26e9723c851c3a1e56b1b1c241d876291a92069086e52774e77890dbc2
size 506
