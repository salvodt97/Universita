version https://git-lfs.github.com/spec/v1
oid sha256:1fd5648bf77752ee2041b5ce5dc25d8b4ca4ed7c2494418d87e0a11257e7e890
size 1134
