version https://git-lfs.github.com/spec/v1
oid sha256:354654b834d035936ba19615a61c72e43bd0a1f9b3f43e7b3168e1bf05a954d8
size 621
