version https://git-lfs.github.com/spec/v1
oid sha256:1206e8895997fb13ca403b48a704ee35cb49f8e0e6d556ea428ce46042b06269
size 851
