version https://git-lfs.github.com/spec/v1
oid sha256:d2c1f23bf0784db5385ca8958d97248df6cf4c77e37e42de0239723b1aa5b85a
size 3076
