version https://git-lfs.github.com/spec/v1
oid sha256:f8d59810ad7a035bcf0863cace1a2de0d57d94c03a5de2d8525d589cc91b4d3d
size 968
