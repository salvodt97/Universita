version https://git-lfs.github.com/spec/v1
oid sha256:cd9bb84ecd786b74cc7e38ee25fdb8106669fafcb15851808fe65c56badf1dab
size 933
