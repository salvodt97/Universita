version https://git-lfs.github.com/spec/v1
oid sha256:ab7e5ef8d5b88c7e3985b041bcdcd1b67339f2be8f31c6ef818164659d3d3dfd
size 5803
