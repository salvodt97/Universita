version https://git-lfs.github.com/spec/v1
oid sha256:11eb565025df414ec466e8136b17780fdabd1ac5ea579738466177d85fadae15
size 727
