version https://git-lfs.github.com/spec/v1
oid sha256:bb65e3eba08d08e76805aa86773c392ef312024da825431a506f4bffcf5bdcf0
size 3464
