version https://git-lfs.github.com/spec/v1
oid sha256:1b0b172938299bce3a9ae8b243b2ceaf34a5cc11c337eb13576f9a8ca60d5327
size 1088
