version https://git-lfs.github.com/spec/v1
oid sha256:f97e8035d4bb030ab83a6138f1d906129111385d508a9fec9fb1736a630778b1
size 444
