version https://git-lfs.github.com/spec/v1
oid sha256:9544f37aaa1248c6ca9ea1081d198c0dc04a48990faa8ce99d653c0e945bf2c3
size 1647
