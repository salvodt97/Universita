version https://git-lfs.github.com/spec/v1
oid sha256:3e33a7f7026e5e5d2c1afc02305452d261b059c37971e7f26bcc85fd89efb2e7
size 1124
