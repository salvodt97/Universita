version https://git-lfs.github.com/spec/v1
oid sha256:b93ba7a2ad1d712cd27d1f760fbd6f42141fd7e4c03fa424d20327351e54fa67
size 1918
