version https://git-lfs.github.com/spec/v1
oid sha256:b5470ac9a41c862a4ebc9b311e9ca9991813141b3d4deea97d014aea18579363
size 887
