version https://git-lfs.github.com/spec/v1
oid sha256:a5db965360e12d319b07c1adf8571212813732b7d5815c318a8259d5802a275e
size 2588
