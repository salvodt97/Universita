version https://git-lfs.github.com/spec/v1
oid sha256:08203f391be3cfe798a19d8bf7d1258f746463f3ce2927fd9dadda6f2975afc8
size 639
