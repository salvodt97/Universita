version https://git-lfs.github.com/spec/v1
oid sha256:2fdec23a9d9ead9caaa90a7beeaa6ab8a014774b3ec035841f30f242ed913c71
size 680
