version https://git-lfs.github.com/spec/v1
oid sha256:3eb89da3e14118e05a33258378ff4fcdd6011176c797a6bae384d3c906610c1c
size 1152
