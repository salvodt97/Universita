version https://git-lfs.github.com/spec/v1
oid sha256:049c3ae1d52a6ae2758dd7d261a4a76c68e9d4ae892b8eb7f3063fc8713f9970
size 2597
