version https://git-lfs.github.com/spec/v1
oid sha256:eb9d28fca128608a8e30f55edff1894058f20f733aaca9a7b4fd062e09c5bdba
size 2105
