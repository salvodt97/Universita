version https://git-lfs.github.com/spec/v1
oid sha256:1ff3410b95f387f7813ad57f65a4c95fbd9ebcd20ca88c5dc233511d747cee64
size 751
