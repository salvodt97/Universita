version https://git-lfs.github.com/spec/v1
oid sha256:7b95a600db52febe8da8e33c0e5b66d30f74717aad8be0b492cd20c730868f9b
size 582
