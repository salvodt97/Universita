version https://git-lfs.github.com/spec/v1
oid sha256:d660e15b2afeeda6d30fd708a125ae7317b9ff78f2235ea0a6048f4c99a88e17
size 3020
