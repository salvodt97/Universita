version https://git-lfs.github.com/spec/v1
oid sha256:9635e34f65096ea6af0e03e725a290af8906d346bb52f912cfa86c24a20fe17a
size 1116
