version https://git-lfs.github.com/spec/v1
oid sha256:d4cf88e20bfec8bf7d7ea98ba22d3d3a20ef08d80e241e41456193d9317097ad
size 1921
