version https://git-lfs.github.com/spec/v1
oid sha256:96b1cc4cb501273da706494a9aac801119a92b5cceada9d89b368a424e1f61f4
size 916
