version https://git-lfs.github.com/spec/v1
oid sha256:cfc6ebf8ab34761f55ac255d3efa35786da3926c26bd24eb8ed9443d4b7bca26
size 4965
