version https://git-lfs.github.com/spec/v1
oid sha256:8702a2294c7ee7f74f1623c2144e15d8ac2de86b717aa6772ea15c16f1dc9ff7
size 1120
