version https://git-lfs.github.com/spec/v1
oid sha256:78045027197100d5adb84ec2646743de7ee903c76737cbeb98ef41054cabf252
size 550
