version https://git-lfs.github.com/spec/v1
oid sha256:72e7715a2fb08d904d82282090082f30373a1ec963fba23c0010ba26fdda06cf
size 1591
