version https://git-lfs.github.com/spec/v1
oid sha256:455263e29bd15b6398a4df6f5f855de136b6b4008b24daf53064a7d3e07e18da
size 1070
