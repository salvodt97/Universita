version https://git-lfs.github.com/spec/v1
oid sha256:a6a7759fcde7bb876e6a59ea9b2e7507cfa9e3e4a5e70a0dc207a294eb166d4f
size 2421
