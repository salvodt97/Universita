version https://git-lfs.github.com/spec/v1
oid sha256:d2682bb9a2ff11ada67fe51c840ac59158c3f9b527ccd9e3d68e8d69574bf144
size 260
