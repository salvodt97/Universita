version https://git-lfs.github.com/spec/v1
oid sha256:fe8277ec25859d71536aa0311ad74603c641394b4b0863d75618c534c439712d
size 382
