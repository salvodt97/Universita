version https://git-lfs.github.com/spec/v1
oid sha256:272a32f56b3fdd9ae063be59e55ada09a524da4b869ab7fe8fd0e6fc43b7ec2c
size 1319
