version https://git-lfs.github.com/spec/v1
oid sha256:675e608006dd9fd6d6e2bc54ae92c72d4eae75721e471b554f8f1c6fa2ad9df4
size 838
