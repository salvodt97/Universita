version https://git-lfs.github.com/spec/v1
oid sha256:b5570c7c9c859ca068f1120df5dad254d095d72d3d00a290878a69687321ca6d
size 1767
