version https://git-lfs.github.com/spec/v1
oid sha256:ae349266c2946029569da972d6729fcb8c1e59675ac90f1f2abf3aa1f965f8f4
size 1183
