version https://git-lfs.github.com/spec/v1
oid sha256:0baf5f61e2360d57e0c20b3794b85a23cd914a0b4a38712098fadf08cf29fdf1
size 271
