version https://git-lfs.github.com/spec/v1
oid sha256:fb9e4208c4fc5a375cacdf465b52aee1fa3a36cb39212841f631dc358b3411f5
size 1239
