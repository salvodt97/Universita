version https://git-lfs.github.com/spec/v1
oid sha256:aa2b6cddc383cf78e309c55f19beb3d30d9d09f479c7c96c3f1f861745146390
size 1854
