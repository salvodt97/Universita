version https://git-lfs.github.com/spec/v1
oid sha256:338832a7dda0b2da008d56d68060a315e9854f80a2de692dee6bd4859ed875e8
size 582
