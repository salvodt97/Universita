version https://git-lfs.github.com/spec/v1
oid sha256:bb7e04813790d9ec43e222f69d8ee2d64f0989000882b3ad52a6a720a67177fb
size 6782
