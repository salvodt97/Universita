version https://git-lfs.github.com/spec/v1
oid sha256:87f8670934401db0b902ad4f409668b803d18508ebc14231c05270bf8a1ff068
size 835
