version https://git-lfs.github.com/spec/v1
oid sha256:08cb5f755c273b8471da31a49b278e0c86f6669328b7124f4438e474795d2ed7
size 789
