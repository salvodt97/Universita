version https://git-lfs.github.com/spec/v1
oid sha256:ee47c52b47df32f06e7cd4de811f6d67b1a0a2c1fc31cc7b5121bb0d9fc0b418
size 262
