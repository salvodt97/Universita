version https://git-lfs.github.com/spec/v1
oid sha256:53f8e2c68792804f276984119744df3195a506f868676f2056396459d18607e4
size 1216
