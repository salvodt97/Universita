version https://git-lfs.github.com/spec/v1
oid sha256:3a2b096fd10e3b070a90c7ba7c310d3a32d2b12547173687914207eb2b7b925c
size 1834
