version https://git-lfs.github.com/spec/v1
oid sha256:3b8f522b01eec591f3b9fe0e8cfce8aae2f0ce30654ec523582e0721ae8a9442
size 897
