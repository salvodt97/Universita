version https://git-lfs.github.com/spec/v1
oid sha256:edd3cfad3f852650e356dc77a84fcae97765dd9ab9e63ab007918d74ffa9d44a
size 3273
