version https://git-lfs.github.com/spec/v1
oid sha256:4692417aa9954e4f235ee707deb7f2533eaaf7b4cae4441d8b7f05e61396e200
size 2205
