version https://git-lfs.github.com/spec/v1
oid sha256:47f066ea622e153d0d5495fbb2d62033446a04e828fa9998bf479b4f9367a311
size 25911
