version https://git-lfs.github.com/spec/v1
oid sha256:851c09f1d8b28cd4499d532e6094a962dd4b0c3b07c999124c9b8fe45a8c621f
size 675
