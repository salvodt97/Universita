version https://git-lfs.github.com/spec/v1
oid sha256:d7306999b3dc082ced9561825906d6717d86bcae1bf67fc754490daf6c3b1244
size 821
