version https://git-lfs.github.com/spec/v1
oid sha256:0b9f29cfa33c26f606e30e0236f7d0ede7f0adc88e93fe1972c4c6b11eed7748
size 1282
