version https://git-lfs.github.com/spec/v1
oid sha256:d560b4c47c26ca524eef559575d1d94aae81f26aeab867af33a7bdbf364e3bfc
size 267
