version https://git-lfs.github.com/spec/v1
oid sha256:855806b56d8a53e70a65e07b215ad2f13222e1e649ba34757af90f58d18fa821
size 324
