version https://git-lfs.github.com/spec/v1
oid sha256:b277fbf1c52c1b47d68621099fde4cd23e14063d5435d4a683f785030057f070
size 459
