version https://git-lfs.github.com/spec/v1
oid sha256:79c497c1bbce6e962d7416708ce466e8deb451fee046c3477b0d06306b2b7098
size 1214
