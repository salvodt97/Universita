version https://git-lfs.github.com/spec/v1
oid sha256:cdf18432a9c57737a69cc11adb27f429fbbc71829c1d10e155b2497f45c1beb9
size 2756
