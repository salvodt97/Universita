version https://git-lfs.github.com/spec/v1
oid sha256:f3845029ae4a7b8d4f99390936fbbadee3d3f89e54c6ea370afb6e91dc0300b0
size 1574
