version https://git-lfs.github.com/spec/v1
oid sha256:4e3914e550d03ca67e0a7bd4bd8d39c7a5675a1ce48293b06912f9914fdab0b4
size 2016
