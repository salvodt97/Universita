version https://git-lfs.github.com/spec/v1
oid sha256:3858fb06e551e4784344f9f97c3068c03c319cec719b8318002235b44c384d95
size 1595
