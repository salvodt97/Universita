version https://git-lfs.github.com/spec/v1
oid sha256:29c96e56c5255af176f818704836c5dcb7c0f99081414778821c020a72e2f5ac
size 715
