version https://git-lfs.github.com/spec/v1
oid sha256:2863b9a1e3a7c4563a323f5284f9343e0a5bd1f2ee887727475d9dbae4bef896
size 1053
