version https://git-lfs.github.com/spec/v1
oid sha256:be6930c37dac5f16b909ebd97943c124aff860ad2036a39c65b9b95a0703529d
size 3221
