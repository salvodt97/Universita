version https://git-lfs.github.com/spec/v1
oid sha256:682c187659fdcf84e59ddec992e0fb8ca8ba868c2e8277fbdd714499c3dd2057
size 498
