version https://git-lfs.github.com/spec/v1
oid sha256:3d645a1def726657ae05f6ea101752bdcb8c27adcb663215038f97f576ea0da6
size 6443
