version https://git-lfs.github.com/spec/v1
oid sha256:7041f05c1f1af07f63e86e85d8f06df26252abfa73646d28a56ac3917d6561c4
size 4120
