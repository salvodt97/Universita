version https://git-lfs.github.com/spec/v1
oid sha256:671c69c3ce4e889fa15cc603df5a38c1555cf060905721b71b2c464d9c3b5b71
size 641
