version https://git-lfs.github.com/spec/v1
oid sha256:54ce62661f295c5ec2d5d92898ed90bee13a68e410e8430628306bffffe78a36
size 935
