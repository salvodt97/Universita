version https://git-lfs.github.com/spec/v1
oid sha256:ea6e2db11d10ed08669a0832a94eb7365f30da1d6118f4d6aec23a0b0372ac78
size 6821
