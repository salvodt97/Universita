version https://git-lfs.github.com/spec/v1
oid sha256:de9d47954ea8b66a5602c65d3e71a3bac1190abd813f2cf35aaff7519a56853c
size 2398
