version https://git-lfs.github.com/spec/v1
oid sha256:e9a2698d7d34465821b01b49fa9c83d2033e956184ae62c568cdf1e9ebc9d23b
size 1130
