version https://git-lfs.github.com/spec/v1
oid sha256:6591d3aad96bbc3db6e796e65ef6949f1302e6c247f4b389edd29666d4950b04
size 1911
