version https://git-lfs.github.com/spec/v1
oid sha256:535c5d4f4b4cd0654ce2f88dc0127614a4b1482072716734102b3b29ceb9fef4
size 3081
