version https://git-lfs.github.com/spec/v1
oid sha256:5407670c18f4bd541a52467997986eae5b0c35bceefcefab6ff949483533cd7f
size 1219
